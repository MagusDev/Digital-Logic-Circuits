

module moore10010(input clk,j,rst,output w);
reg [2:0]ns;
reg [2:0]ps;

parameter [2:0]A=3'b000,B=3'b001,C=3'b010,D=3'b011,E=3'b100, F=3'b101;

always @(ps,j) begin


case(ps)
A: ns = j? B : A;
B: ns = j? B : C;
C: ns = j? B : D;
D: ns = j? E : A;
E: ns = j? B : F;
F: ns = j? B : D;
default: ns =A;
 endcase
end 

assign w = (ps == F) ? 1'b1 : 1'b0;
always @(posedge clk,posedge rst) begin

if (rst)
ps<= 3'b000;
else
ps<= ns;
end

endmodule
